library ieee;
use ieee.std_logic_1164.all;

ENTITY EVEN_DETECTOR_TESTBENCH is
end EVEN_DETECTOR_TESTBENCH;

architecture TB_ARCH OF EVEN_DETECTOR_TESTBENCH is
	component EVEN_DETECTOR_TESTBENCH
		PORT(
			A: IN STD_LOGIC_VECTOR(2 downto 0);
			EVEN: OUT std_logic_1164
		);
	END component;
	SIGNAL TEST_IN : STD_LOGIC_VECTOR(2 downto0);
	SIGNAL TEST_OUT: STD_LOGIC;
	
BEGIN
	-- INSTATNTIATE THE CIRCUIT UNDER TEST 
	UUT: EVEN_DETECTOR 
		PORT MAP(A=>TEST_IN, EVEN => TEST_OUT);
	-- TEST VECTOR GENERATOR
	process
	BEGIN
		TEST_IN	<= "000";
		WAIT FOR 200 ns;
		TEST_IN	<= "001";
		WAIT FOR 200 ns;
		TEST_IN	<= "010";
		WAIT FOR 200 ns;
		TEST_IN	<= "011";
		WAIT FOR 200 ns;
		TEST_IN	<= "100";
		WAIT FOR 200 ns;
		TEST_IN	<= "101";
		WAIT FOR 200 ns;
		TEST_IN	<= "110";
		WAIT FOR 200 ns;
		TEST_IN	<= "111";
		WAIT FOR 200 ns;
	END PROCESS;
	-- VERIFIER
	PROCESS
		VARIABLE ERROR_STATUS : BOOLEAN;
	BEGIN
		WAIT ON TEST_IN;
		WAIT FOR 100 ns;
		IF ((TEST_IN = "000" AND TEST_OUT='1') OR
			(TEST_IN = "001" AND TEST_OUT='0') OR
			(TEST_IN = "010" AND TEST_OUT='0') OR
			(TEST_IN = "011" AND TEST_OUT='1') OR
			(TEST_IN = "100" AND TEST_OUT='0') OR
			(TEST_IN = "101" AND TEST_OUT='1') OR
			(TEST_IN = "110" AND TEST_OUT='1') OR
			(TEST_IN = "111" AND TEST_OUT='0'))
		THEN 
			ERROR_STATUS := FALSE;
		ELSE 
			ERROR_STATUS := TRUE;
		END IF;
		-- ERROR REPORTING
		ASSERT NOT ERROR_STATUS
			REPORT "TEST FAILED."
			SEVERITY NOTE;
	END PROCESS;
END TB_ARCH;
